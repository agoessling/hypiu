`ifndef ALU_CODE_H_
`define ALU_CODE_H_

`define ALU_BIT_NUM 4

`define ALU_ZERO    0
`define ALU_A       1
`define ALU_B       2
`define ALU_ADD     3
`define ALU_SUB     4

`endif
