`ifndef OPCODE_VH_
`define OPCODE_VH_

`define OPCODE_LDI   0
`define OPCODE_STI   1
`define OPCODE_ADD   2
`define OPCODE_SUB   3
`define OPCODE_ADDI  4
`define OPCODE_SUBI  5
`define OPCODE_MOV   6
`define OPCODE_BRZ   7
`define OPCODE_JMP   8

`endif
